/*
 *  addr_gen.sv -- address generator for multi-bank memories incl. registers
 *  ETRI <SW-SoC AI Deep Learning HW Accelerator RTL Design> course material
 *
 *  first draft by Junyoung Park
 */

`timescale 1ns / 1ps

module addr_gen #(
  parameter integer ADDR_WIDTH = 12,
  parameter integer DATA_WIDTH = 32
  ) (
  // clock and resetn from domain a
  input  wire clk_a,
  input  wire arstz_aq,

  // signals from the external interfaces
  cnnip_mem_if.slave  from_axi4l_mem_if,

  // signals to the internal interfaces
  cnnip_mem_if.master to_register_if,
  cnnip_mem_if.master to_input_mem_if,
  cnnip_mem_if.master to_weight_mem_if,
  cnnip_mem_if.master to_feature_mem_if
  );

  wire to_register;
  wire to_input_mem;
  wire to_weight_mem;
  wire to_feature_mem;

  wire [3:0] select;

  // address multiplexer
  assign to_register    = (from_axi4l_mem_if.addr[11:8] == 4'h0) ? 1: 0;
  assign to_input_mem   = (from_axi4l_mem_if.addr[11:8] == 4'h1) ? 1: 0;
  assign to_weight_mem  = (from_axi4l_mem_if.addr[11:8] == 4'h2) ? 1: 0;
  assign to_feature_mem = (from_axi4l_mem_if.addr[11:8] == 4'h3) ? 1: 0;

  assign select = { to_feature_mem,
                    to_weight_mem,
                    to_input_mem,
                    to_register };

  assign to_register_if.en   = (to_register == 1) ? from_axi4l_mem_if.en   : 'b0;
  assign to_register_if.we   = (to_register == 1) ? from_axi4l_mem_if.we   : 'b0;
  assign to_register_if.addr = (to_register == 1) ? from_axi4l_mem_if.addr : 'b0;
  assign to_register_if.din  = (to_register == 1) ? from_axi4l_mem_if.din  : 'b0;

  assign to_input_mem_if.en   = (to_input_mem == 1) ? from_axi4l_mem_if.en   : 'b0;
  assign to_input_mem_if.we   = (to_input_mem == 1) ? from_axi4l_mem_if.we   : 'b0;
  assign to_input_mem_if.addr = (to_input_mem == 1) ? from_axi4l_mem_if.addr : 'b0;
  assign to_input_mem_if.din  = (to_input_mem == 1) ? from_axi4l_mem_if.din  : 'b0;

  assign to_weight_mem_if.en   = (to_weight_mem == 1) ? from_axi4l_mem_if.en   : 'b0;
  assign to_weight_mem_if.we   = (to_weight_mem == 1) ? from_axi4l_mem_if.we   : 'b0;
  assign to_weight_mem_if.addr = (to_weight_mem == 1) ? from_axi4l_mem_if.addr : 'b0;
  assign to_weight_mem_if.din  = (to_weight_mem == 1) ? from_axi4l_mem_if.din  : 'b0;

  assign to_feature_mem_if.en   = (to_feature_mem == 1) ? from_axi4l_mem_if.en   : 'b0;
  assign to_feature_mem_if.we   = (to_feature_mem == 1) ? from_axi4l_mem_if.we   : 'b0;
  assign to_feature_mem_if.addr = (to_feature_mem == 1) ? from_axi4l_mem_if.addr : 'b0;
  assign to_feature_mem_if.din  = (to_feature_mem == 1) ? from_axi4l_mem_if.din  : 'b0;
/*
  assign from_axi4l_mem_if.dout = (to_register == 1) ? to_register_if.dout :
                                  (to_input_mem == 1) ? to_input_mem_if.dout :
                                  (to_weight_mem == 1) ? to_weight_mem_if.dout :
                                  (to_feature_mem == 1) ? to_feature_mem_if.dout : 0;
                                  
  assign from_axi4l_mem_if.valid = (to_register == 1) ? to_register_if.valid :
                                   (to_input_mem == 1) ? to_input_mem_if.valid :
                                   (to_weight_mem == 1) ? to_weight_mem_if.valid :
                                   (to_feature_mem == 1) ? to_feature_mem_if.valid : 0;
*/
//always_comb
//begin
//    if(to_register == 1)
//        from_axi4l_mem_if.dout = to_register_if.dout;
//    else if(to_input_mem == 1)
//        from_axi4l_mem_if.dout = to_input_mem_if.dout;
//    else if(to_weight_mem == 1)
//        from_axi4l_mem_if.dout = to_weight_mem_if.dout;
//    else if(to_feature_mem == 1)
//        from_axi4l_mem_if.dout = to_feature_mem_if.dout;
//    else
//        from_axi4l_mem_if.dout = 0;
//end
//always_comb
//begin
//    if(to_register == 1)
//        from_axi4l_mem_if.valid = to_register_if.valid;
//    else if(to_input_mem == 1)
//        from_axi4l_mem_if.valid = to_input_mem_if.valid;
//    else if(to_weight_mem == 1)
//        from_axi4l_mem_if.valid = to_weight_mem_if.valid;
//    else if(to_feature_mem == 1)
//        from_axi4l_mem_if.valid = to_feature_mem_if.valid;
//    else
//        from_axi4l_mem_if.valid = 0;
//end


  always_comb // always @(*)
  begin
    // unfortunately, the current vivado does not support unique case syntax
    // unique case(select)
    from_axi4l_mem_if.dout = 0;
    case(select)
              // 0: from_axi4l_mem_if.dout = 0;
      4'b0001: from_axi4l_mem_if.dout = to_register_if.dout;
      4'b0010: from_axi4l_mem_if.dout = to_input_mem_if.dout;
      4'b0100: from_axi4l_mem_if.dout = to_weight_mem_if.dout;
      4'b1000: from_axi4l_mem_if.dout = to_feature_mem_if.dout;
      // {4{1'bx}}: from_axi4l_mem_if.dout = 0;
    endcase
  end

  always_comb
  begin
    // unique case(select)
    from_axi4l_mem_if.valid = 0;
    case(select)
              // 0: from_axi4l_mem_if.valid = 0;
      4'b0001: from_axi4l_mem_if.valid = to_register_if.valid;
      4'b0010: from_axi4l_mem_if.valid = to_input_mem_if.valid;
      4'b0100: from_axi4l_mem_if.valid = to_weight_mem_if.valid;
      4'b1000: from_axi4l_mem_if.valid = to_feature_mem_if.valid;
      // {4{1'bx}}: from_axi4l_mem_if.valid = 0;
    endcase
  end

endmodule
